// avalon_jtag.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module avalon_jtag (
		output wire [16:0] AVL_MM_slave_0_avs_s0_address,     // AVL_MM_slave_0_avs_s0.address
		output wire        AVL_MM_slave_0_avs_s0_read,        //                      .read
		input  wire [7:0]  AVL_MM_slave_0_avs_s0_readdata,    //                      .readdata
		output wire        AVL_MM_slave_0_avs_s0_write,       //                      .write
		output wire [7:0]  AVL_MM_slave_0_avs_s0_writedata,   //                      .writedata
		input  wire        AVL_MM_slave_0_avs_s0_waitrequest, //                      .waitrequest
		output wire        AVL_MM_slave_0_reset_reset,        //  AVL_MM_slave_0_reset.reset
		input  wire        clk_clk,                           //                   clk.clk
		input  wire        reset_reset_n                      //                 reset.reset_n
	);

	wire  [31:0] master_0_master_readdata;      // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;   // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;       // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire         master_0_master_read;          // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire   [3:0] master_0_master_byteenable;    // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire         master_0_master_readdatavalid; // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;         // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire  [31:0] master_0_master_writedata;     // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata

	avalon_jtag_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_clk),                       //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                //    clk_reset.reset
		.master_address       (master_0_master_address),       //       master.address
		.master_readdata      (master_0_master_readdata),      //             .readdata
		.master_read          (master_0_master_read),          //             .read
		.master_write         (master_0_master_write),         //             .write
		.master_writedata     (master_0_master_writedata),     //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                               // master_reset.reset
	);

	avalon_jtag_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                           //                                  clk_0_clk.clk
		.AVL_MM_slave_0_reset_reset_bridge_in_reset_reset (AVL_MM_slave_0_reset_reset),        // AVL_MM_slave_0_reset_reset_bridge_in_reset.reset
		.master_0_clk_reset_reset_bridge_in_reset_reset   (AVL_MM_slave_0_reset_reset),        //   master_0_clk_reset_reset_bridge_in_reset.reset
		.master_0_master_address                          (master_0_master_address),           //                            master_0_master.address
		.master_0_master_waitrequest                      (master_0_master_waitrequest),       //                                           .waitrequest
		.master_0_master_byteenable                       (master_0_master_byteenable),        //                                           .byteenable
		.master_0_master_read                             (master_0_master_read),              //                                           .read
		.master_0_master_readdata                         (master_0_master_readdata),          //                                           .readdata
		.master_0_master_readdatavalid                    (master_0_master_readdatavalid),     //                                           .readdatavalid
		.master_0_master_write                            (master_0_master_write),             //                                           .write
		.master_0_master_writedata                        (master_0_master_writedata),         //                                           .writedata
		.AVL_MM_slave_0_avs_s0_address                    (AVL_MM_slave_0_avs_s0_address),     //                      AVL_MM_slave_0_avs_s0.address
		.AVL_MM_slave_0_avs_s0_write                      (AVL_MM_slave_0_avs_s0_write),       //                                           .write
		.AVL_MM_slave_0_avs_s0_read                       (AVL_MM_slave_0_avs_s0_read),        //                                           .read
		.AVL_MM_slave_0_avs_s0_readdata                   (AVL_MM_slave_0_avs_s0_readdata),    //                                           .readdata
		.AVL_MM_slave_0_avs_s0_writedata                  (AVL_MM_slave_0_avs_s0_writedata),   //                                           .writedata
		.AVL_MM_slave_0_avs_s0_waitrequest                (AVL_MM_slave_0_avs_s0_waitrequest)  //                                           .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),             // reset_in0.reset
		.clk            (clk_clk),                    //       clk.clk
		.reset_out      (AVL_MM_slave_0_reset_reset), // reset_out.reset
		.reset_req      (),                           // (terminated)
		.reset_req_in0  (1'b0),                       // (terminated)
		.reset_in1      (1'b0),                       // (terminated)
		.reset_req_in1  (1'b0),                       // (terminated)
		.reset_in2      (1'b0),                       // (terminated)
		.reset_req_in2  (1'b0),                       // (terminated)
		.reset_in3      (1'b0),                       // (terminated)
		.reset_req_in3  (1'b0),                       // (terminated)
		.reset_in4      (1'b0),                       // (terminated)
		.reset_req_in4  (1'b0),                       // (terminated)
		.reset_in5      (1'b0),                       // (terminated)
		.reset_req_in5  (1'b0),                       // (terminated)
		.reset_in6      (1'b0),                       // (terminated)
		.reset_req_in6  (1'b0),                       // (terminated)
		.reset_in7      (1'b0),                       // (terminated)
		.reset_req_in7  (1'b0),                       // (terminated)
		.reset_in8      (1'b0),                       // (terminated)
		.reset_req_in8  (1'b0),                       // (terminated)
		.reset_in9      (1'b0),                       // (terminated)
		.reset_req_in9  (1'b0),                       // (terminated)
		.reset_in10     (1'b0),                       // (terminated)
		.reset_req_in10 (1'b0),                       // (terminated)
		.reset_in11     (1'b0),                       // (terminated)
		.reset_req_in11 (1'b0),                       // (terminated)
		.reset_in12     (1'b0),                       // (terminated)
		.reset_req_in12 (1'b0),                       // (terminated)
		.reset_in13     (1'b0),                       // (terminated)
		.reset_req_in13 (1'b0),                       // (terminated)
		.reset_in14     (1'b0),                       // (terminated)
		.reset_req_in14 (1'b0),                       // (terminated)
		.reset_in15     (1'b0),                       // (terminated)
		.reset_req_in15 (1'b0)                        // (terminated)
	);

endmodule
